module cordic_floatingpoint_mul_K_Left_shifter (
	//	Inputs
	input	[47:0]	in,
	input	[4:0]	shift,
	
	//	Output
	output	[22:0]	out
);

/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
 
 //	Stage 1 <<16
 wire	[37:0]	stage1;
 
 //	Stage 2 <<8
 wire	[29:0]	stage2;
 
 //	Stage 3 <<4
 wire	[25:0]	stage3;
 
 //	Stage 4 <<2
 wire	[23:0]	stage4;
 
 //	Stage 5 <<1
 wire	[22:0]	stage5;
 
/*****************************************************************************
 *                            Stage 1 shift 16                               *
 *****************************************************************************/
 
 assign stage1[37:7] = (shift[4]) ? in[30:0] : in[46:16];
 assign stage1[6] = !shift[4] & in[15];
 assign stage1[5] = !shift[4] & in[14];
 assign stage1[4] = !shift[4] & in[13];
 assign stage1[3] = !shift[4] & in[12];
 assign stage1[2] = !shift[4] & in[11];
 assign stage1[1] = !shift[4] & in[10];
 assign stage1[0] = !shift[4] & in[9];
 
/*****************************************************************************
 *                            Stage 2 shift 8                                *
 *****************************************************************************/
 
 assign stage2 = (shift[3]) ? stage1[29:0] : stage1[37:8];
 
/*****************************************************************************
 *                            Stage 3 shift 4                                *
 *****************************************************************************/
 
 assign stage3 = (shift[2]) ? stage2[25:0] : stage2[29:4];
 
/*****************************************************************************
 *                            Stage 4 shift 2                                *
 *****************************************************************************/
 
 assign stage4 = (shift[1]) ? stage3[23:0] : stage3[25:2];
 
/*****************************************************************************
 *                            Stage 5 shift 1                                *
 *****************************************************************************/
 
 assign stage5 = (shift[0]) ? stage4[22:0] : stage4[23:1];
 
 assign out = stage5;
 
endmodule
